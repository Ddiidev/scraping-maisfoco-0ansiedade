module models

pub type ThumbLink = string
