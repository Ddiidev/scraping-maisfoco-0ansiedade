module models

pub enum MultimediaMode {
	search_tv
	search_movie
}
