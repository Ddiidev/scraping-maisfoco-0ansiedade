module wcontext

import veb

pub struct WsCtx {
	veb.Context
}
