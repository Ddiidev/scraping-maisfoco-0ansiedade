module components

import slices.shareds.components.badge

pub struct Components {
	badge.Badge
}