module models

pub type TrailerLink = string
